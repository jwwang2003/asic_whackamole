// defines.vh
`ifndef DEFINES_VH
`define DEFINES_VH

// … other macros …

//-----------------------------------------------------------------------------
// Define a 50 kHz clock frequency (in Hertz)
//-----------------------------------------------------------------------------
`define CLK_FREQ 50_000

`endif
